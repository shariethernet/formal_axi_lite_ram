bind axil_ram f_axil inst_1(
          clk,
          rst,
      s_axil_awaddr,
          s_axil_awprot,
          s_axil_awvalid,
         s_axil_awready,
  s_axil_wdata,
          s_axil_wstrb,
          s_axil_wvalid,
         s_axil_wready,
 s_axil_bresp,
         s_axil_bvalid,
          s_axil_bready,
  s_axil_araddr,
          s_axil_arprot,
          s_axil_arvalid,
         s_axil_arready,
 s_axil_rdata,
         s_axil_rresp,
         s_axil_rvalid,
          s_axil_rready
);